library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity BLDCCtrl is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity;

architecture rtl of BLDCCtrl is

begin

    

end architecture;